library verilog;
use verilog.vl_types.all;
entity UpDownCounter_8bitExample_vlg_vec_tst is
end UpDownCounter_8bitExample_vlg_vec_tst;
