library verilog;
use verilog.vl_types.all;
entity UpDownCounter_8bit_tb is
end UpDownCounter_8bit_tb;
