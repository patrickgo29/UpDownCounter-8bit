library verilog;
use verilog.vl_types.all;
entity UpDownCounter_8bit_vlg_vec_tst is
end UpDownCounter_8bit_vlg_vec_tst;
